`timescale 1ns / 1ps

module DB(input[31:0] in,output reg [31:0] out);


		reg [7:0] exp;
		reg sign;
		reg [22:0]frac;
		
		reg[1:0]  in_status ;
		
	   localparam usual = 2'b00;
	   localparam zero = 2'b01;
	   localparam inf = 2'b10;
	   localparam nan = 2'b11;
		

		
		reg res_sgn;
		reg [7:0]  res_exp;
		reg [22:0] res_frac;
		
		reg [31:0] log1f;
		reg [31:0] exp_formatted;  //(e-127)*log2
		wire [31:0] tmp_res;

		ADD A0 (.opr1(log1f),.opr2(exp_formatted),.res(tmp_res));
always @(*) begin

    sign = in[31] ;
    exp = in[30:23];
    frac = in[22:0] ;
	 
		case (frac[22:18])
            0: log1f = 32'b00000000000000000000000000000000;
            1: log1f = 32'b00111110100010001101100011010010;
            2: log1f = 32'b00111111000001101100110111011110;
            3: log1f = 32'b00111111010001110100001010110000;
            4: log1f = 32'b00111111100000101111001101010001;
            5: log1f = 32'b00111111101000010110100110011000;
            6: log1f = 32'b00111111101111110000111111100100;
            7: log1f = 32'b00111111110110111111000100000010;
            8: log1f = 32'b00111111111110000001011011110010;
            9: log1f = 32'b01000000000010011100010101111000;
            10: log1f = 32'b01000000000101110010101011001000;
            11: log1f = 32'b01000000001001000011111101100110;
            12: log1f = 32'b01000000001100010000011100000111;
            13: log1f = 32'b01000000001111011000010100100010;
            14: log1f = 32'b01000000010010011011110011110001;
            15: log1f = 32'b01000000010101011011000101111100;
            16: log1f = 32'b01000000011000010110010110010101;
            17: log1f = 32'b01000000011011001101101111101000;
            18: log1f = 32'b01000000011110000001011011110010;
            19: log1f = 32'b01000000100000011000110010000111;
            20: log1f = 32'b01000000100001101111001000110111;
            21: log1f = 32'b01000000100011000011110110010110;
            22: log1f = 32'b01000000100100010110111110011111;
            23: log1f = 32'b01000000100101101000100101000000;
            24: log1f = 32'b01000000100110111000101101011010;
            25: log1f = 32'b01000000101000000111011011000100;
            26: log1f = 32'b01000000101001010100110001000101;
            27: log1f = 32'b01000000101010100000110010011111;
            28: log1f = 32'b01000000101011101011100010001000;
            29: log1f = 32'b01000000101100110101000010101011;
            30: log1f = 32'b01000000101101111101010110101110;
            31: log1f = 32'b01000000101111000100100000110000;
        endcase
		
		case(exp)
		    0: log1f = 32'b11000100001111110010011101110000;
        1: log1f = 32'b11000100001111011010011000011110;
        2: log1f = 32'b11000100001111000010010011001101;
        3: log1f = 32'b11000100001110101010001101111011;
        4: log1f = 32'b11000100001110010010001000101010;
        5: log1f = 32'b11000100001101111010000011011000;
        6: log1f = 32'b11000100001101100001111110000111;
        7: log1f = 32'b11000100001101001001111000110101;
        8: log1f = 32'b11000100001100110001110011100100;
        9: log1f = 32'b11000100001100011001101110010010;
        10: log1f = 32'b11000100001100000001101001000001;
        11: log1f = 32'b11000100001011101001100011101111;
        12: log1f = 32'b11000100001011010001011110011110;
        13: log1f = 32'b11000100001010111001011001001100;
        14: log1f = 32'b11000100001010100001010011111011;
        15: log1f = 32'b11000100001010001001001110101001;
        16: log1f = 32'b11000100001001110001001001010111;
        17: log1f = 32'b11000100001001011001000100000110;
        18: log1f = 32'b11000100001001000000111110110100;
        19: log1f = 32'b11000100001000101000111001100011;
        20: log1f = 32'b11000100001000010000110100010001;
        21: log1f = 32'b11000100000111111000101111000000;
        22: log1f = 32'b11000100000111100000101001101110;
        23: log1f = 32'b11000100000111001000100100011101;
        24: log1f = 32'b11000100000110110000011111001011;
        25: log1f = 32'b11000100000110011000011001111010;
        26: log1f = 32'b11000100000110000000010100101000;
        27: log1f = 32'b11000100000101101000001111010111;
        28: log1f = 32'b11000100000101010000001010000101;
        29: log1f = 32'b11000100000100111000000100110100;
        30: log1f = 32'b11000100000100011111111111100010;
        31: log1f = 32'b11000100000100000111111010010001;
        32: log1f = 32'b11000100000011101111110100111111;
        33: log1f = 32'b11000100000011010111101111101110;
        34: log1f = 32'b11000100000010111111101010011100;
        35: log1f = 32'b11000100000010100111100101001011;
        36: log1f = 32'b11000100000010001111011111111001;
        37: log1f = 32'b11000100000001110111011010101000;
        38: log1f = 32'b11000100000001011111010101010110;
        39: log1f = 32'b11000100000001000111010000000101;
        40: log1f = 32'b11000100000000101111001010110011;
        41: log1f = 32'b11000100000000010111000101100010;
        42: log1f = 32'b11000011111111111110000000100001;
        43: log1f = 32'b11000011111111001101110101111110;
        44: log1f = 32'b11000011111110011101101011011010;
        45: log1f = 32'b11000011111101101101100000110111;
        46: log1f = 32'b11000011111100111101010110010100;
        47: log1f = 32'b11000011111100001101001011110001;
        48: log1f = 32'b11000011111011011101000001001110;
        49: log1f = 32'b11000011111010101100110110101011;
        50: log1f = 32'b11000011111001111100101100001000;
        51: log1f = 32'b11000011111001001100100001100101;
        52: log1f = 32'b11000011111000011100010111000010;
        53: log1f = 32'b11000011110111101100001100011111;
        54: log1f = 32'b11000011110110111100000001111100;
        55: log1f = 32'b11000011110110001011110111011001;
        56: log1f = 32'b11000011110101011011101100110110;
        57: log1f = 32'b11000011110100101011100010010011;
        58: log1f = 32'b11000011110011111011010111110000;
        59: log1f = 32'b11000011110011001011001101001101;
        60: log1f = 32'b11000011110010011011000010101010;
        61: log1f = 32'b11000011110001101010111000000111;
        62: log1f = 32'b11000011110000111010101101100100;
        63: log1f = 32'b11000011110000001010100011000001;
        64: log1f = 32'b11000011101111011010011000011110;
        65: log1f = 32'b11000011101110101010001101111011;
        66: log1f = 32'b11000011101101111010000011011000;
        67: log1f = 32'b11000011101101001001111000110101;
        68: log1f = 32'b11000011101100011001101110010010;
        69: log1f = 32'b11000011101011101001100011101111;
        70: log1f = 32'b11000011101010111001011001001100;
        71: log1f = 32'b11000011101010001001001110101001;
        72: log1f = 32'b11000011101001011001000100000110;
        73: log1f = 32'b11000011101000101000111001100011;
        74: log1f = 32'b11000011100111111000101111000000;
        75: log1f = 32'b11000011100111001000100100011101;
        76: log1f = 32'b11000011100110011000011001111010;
        77: log1f = 32'b11000011100101101000001111010111;
        78: log1f = 32'b11000011100100111000000100110100;
        79: log1f = 32'b11000011100100000111111010010001;
        80: log1f = 32'b11000011100011010111101111101110;
        81: log1f = 32'b11000011100010100111100101001011;
        82: log1f = 32'b11000011100001110111011010101000;
        83: log1f = 32'b11000011100001000111010000000101;
        84: log1f = 32'b11000011100000010111000101100010;
        85: log1f = 32'b11000011011111001101110101111110;
        86: log1f = 32'b11000011011101101101100000110111;
        87: log1f = 32'b11000011011100001101001011110001;
        88: log1f = 32'b11000011011010101100110110101011;
        89: log1f = 32'b11000011011001001100100001100101;
        90: log1f = 32'b11000011010111101100001100011111;
        91: log1f = 32'b11000011010110001011110111011001;
        92: log1f = 32'b11000011010100101011100010010011;
        93: log1f = 32'b11000011010011001011001101001101;
        94: log1f = 32'b11000011010001101010111000000111;
        95: log1f = 32'b11000011010000001010100011000001;
        96: log1f = 32'b11000011001110101010001101111011;
        97: log1f = 32'b11000011001101001001111000110101;
        98: log1f = 32'b11000011001011101001100011101111;
        99: log1f = 32'b11000011001010001001001110101001;
        100: log1f = 32'b11000011001000101000111001100011;
        101: log1f = 32'b11000011000111001000100100011101;
        102: log1f = 32'b11000011000101101000001111010111;
        103: log1f = 32'b11000011000100000111111010010001;
        104: log1f = 32'b11000011000010100111100101001011;
        105: log1f = 32'b11000011000001000111010000000101;
        106: log1f = 32'b11000010111111001101110101111110;
        107: log1f = 32'b11000010111100001101001011110001;
        108: log1f = 32'b11000010111001001100100001100101;
        109: log1f = 32'b11000010110110001011110111011001;
        110: log1f = 32'b11000010110011001011001101001101;
        111: log1f = 32'b11000010110000001010100011000001;
        112: log1f = 32'b11000010101101001001111000110101;
        113: log1f = 32'b11000010101010001001001110101001;
        114: log1f = 32'b11000010100111001000100100011101;
        115: log1f = 32'b11000010100100000111111010010001;
        116: log1f = 32'b11000010100001000111010000000101;
        117: log1f = 32'b11000010011100001101001011110001;
        118: log1f = 32'b11000010010110001011110111011001;
        119: log1f = 32'b11000010010000001010100011000001;
        120: log1f = 32'b11000010001010001001001110101001;
        121: log1f = 32'b11000010000100000111111010010001;
        122: log1f = 32'b11000001111100001101001011110001;
        123: log1f = 32'b11000001110000001010100011000001;
        124: log1f = 32'b11000001100100000111111010010001;
        125: log1f = 32'b11000001010000001010100011000001;
        126: log1f = 32'b11000000110000001010100011000001;
        127: log1f = 32'b00000000000000000000000000000000;
        128: log1f = 32'b01000000110000001010100011000001;
        129: log1f = 32'b01000001010000001010100011000001;
        130: log1f = 32'b01000001100100000111111010010001;
        131: log1f = 32'b01000001110000001010100011000001;
        132: log1f = 32'b01000001111100001101001011110001;
        133: log1f = 32'b01000010000100000111111010010001;
        134: log1f = 32'b01000010001010001001001110101001;
        135: log1f = 32'b01000010010000001010100011000001;
        136: log1f = 32'b01000010010110001011110111011001;
        137: log1f = 32'b01000010011100001101001011110001;
        138: log1f = 32'b01000010100001000111010000000101;
        139: log1f = 32'b01000010100100000111111010010001;
        140: log1f = 32'b01000010100111001000100100011101;
        141: log1f = 32'b01000010101010001001001110101001;
        142: log1f = 32'b01000010101101001001111000110101;
        143: log1f = 32'b01000010110000001010100011000001;
        144: log1f = 32'b01000010110011001011001101001101;
        145: log1f = 32'b01000010110110001011110111011001;
        146: log1f = 32'b01000010111001001100100001100101;
        147: log1f = 32'b01000010111100001101001011110001;
        148: log1f = 32'b01000010111111001101110101111110;
        149: log1f = 32'b01000011000001000111010000000101;
        150: log1f = 32'b01000011000010100111100101001011;
        151: log1f = 32'b01000011000100000111111010010001;
        152: log1f = 32'b01000011000101101000001111010111;
        153: log1f = 32'b01000011000111001000100100011101;
        154: log1f = 32'b01000011001000101000111001100011;
        155: log1f = 32'b01000011001010001001001110101001;
        156: log1f = 32'b01000011001011101001100011101111;
        157: log1f = 32'b01000011001101001001111000110101;
        158: log1f = 32'b01000011001110101010001101111011;
        159: log1f = 32'b01000011010000001010100011000001;
        160: log1f = 32'b01000011010001101010111000000111;
        161: log1f = 32'b01000011010011001011001101001101;
        162: log1f = 32'b01000011010100101011100010010011;
        163: log1f = 32'b01000011010110001011110111011001;
        164: log1f = 32'b01000011010111101100001100011111;
        165: log1f = 32'b01000011011001001100100001100101;
        166: log1f = 32'b01000011011010101100110110101011;
        167: log1f = 32'b01000011011100001101001011110001;
        168: log1f = 32'b01000011011101101101100000110111;
        169: log1f = 32'b01000011011111001101110101111110;
        170: log1f = 32'b01000011100000010111000101100010;
        171: log1f = 32'b01000011100001000111010000000101;
        172: log1f = 32'b01000011100001110111011010101000;
        173: log1f = 32'b01000011100010100111100101001011;
        174: log1f = 32'b01000011100011010111101111101110;
        175: log1f = 32'b01000011100100000111111010010001;
        176: log1f = 32'b01000011100100111000000100110100;
        177: log1f = 32'b01000011100101101000001111010111;
        178: log1f = 32'b01000011100110011000011001111010;
        179: log1f = 32'b01000011100111001000100100011101;
        180: log1f = 32'b01000011100111111000101111000000;
        181: log1f = 32'b01000011101000101000111001100011;
        182: log1f = 32'b01000011101001011001000100000110;
        183: log1f = 32'b01000011101010001001001110101001;
        184: log1f = 32'b01000011101010111001011001001100;
        185: log1f = 32'b01000011101011101001100011101111;
        186: log1f = 32'b01000011101100011001101110010010;
        187: log1f = 32'b01000011101101001001111000110101;
        188: log1f = 32'b01000011101101111010000011011000;
        189: log1f = 32'b01000011101110101010001101111011;
        190: log1f = 32'b01000011101111011010011000011110;
        191: log1f = 32'b01000011110000001010100011000001;
        192: log1f = 32'b01000011110000111010101101100100;
        193: log1f = 32'b01000011110001101010111000000111;
        194: log1f = 32'b01000011110010011011000010101010;
        195: log1f = 32'b01000011110011001011001101001101;
        196: log1f = 32'b01000011110011111011010111110000;
        197: log1f = 32'b01000011110100101011100010010011;
        198: log1f = 32'b01000011110101011011101100110110;
        199: log1f = 32'b01000011110110001011110111011001;
        200: log1f = 32'b01000011110110111100000001111100;
        201: log1f = 32'b01000011110111101100001100011111;
        202: log1f = 32'b01000011111000011100010111000010;
        203: log1f = 32'b01000011111001001100100001100101;
        204: log1f = 32'b01000011111001111100101100001000;
        205: log1f = 32'b01000011111010101100110110101011;
        206: log1f = 32'b01000011111011011101000001001110;
        207: log1f = 32'b01000011111100001101001011110001;
        208: log1f = 32'b01000011111100111101010110010100;
        209: log1f = 32'b01000011111101101101100000110111;
        210: log1f = 32'b01000011111110011101101011011010;
        211: log1f = 32'b01000011111111001101110101111110;
        212: log1f = 32'b01000011111111111110000000100001;
        213: log1f = 32'b01000100000000010111000101100010;
        214: log1f = 32'b01000100000000101111001010110011;
        215: log1f = 32'b01000100000001000111010000000101;
        216: log1f = 32'b01000100000001011111010101010110;
        217: log1f = 32'b01000100000001110111011010101000;
        218: log1f = 32'b01000100000010001111011111111001;
        219: log1f = 32'b01000100000010100111100101001011;
        220: log1f = 32'b01000100000010111111101010011100;
        221: log1f = 32'b01000100000011010111101111101110;
        222: log1f = 32'b01000100000011101111110100111111;
        223: log1f = 32'b01000100000100000111111010010001;
        224: log1f = 32'b01000100000100011111111111100010;
        225: log1f = 32'b01000100000100111000000100110100;
        226: log1f = 32'b01000100000101010000001010000101;
        227: log1f = 32'b01000100000101101000001111010111;
        228: log1f = 32'b01000100000110000000010100101000;
        229: log1f = 32'b01000100000110011000011001111010;
        230: log1f = 32'b01000100000110110000011111001011;
        231: log1f = 32'b01000100000111001000100100011101;
        232: log1f = 32'b01000100000111100000101001101110;
        233: log1f = 32'b01000100000111111000101111000000;
        234: log1f = 32'b01000100001000010000110100010001;
        235: log1f = 32'b01000100001000101000111001100011;
        236: log1f = 32'b01000100001001000000111110110100;
        237: log1f = 32'b01000100001001011001000100000110;
        238: log1f = 32'b01000100001001110001001001010111;
        239: log1f = 32'b01000100001010001001001110101001;
        240: log1f = 32'b01000100001010100001010011111011;
        241: log1f = 32'b01000100001010111001011001001100;
        242: log1f = 32'b01000100001011010001011110011110;
        243: log1f = 32'b01000100001011101001100011101111;
        244: log1f = 32'b01000100001100000001101001000001;
        245: log1f = 32'b01000100001100011001101110010010;
        246: log1f = 32'b01000100001100110001110011100100;
        247: log1f = 32'b01000100001101001001111000110101;
        248: log1f = 32'b01000100001101100001111110000111;
        249: log1f = 32'b01000100001101111010000011011000;
        250: log1f = 32'b01000100001110010010001000101010;
        251: log1f = 32'b01000100001110101010001101111011;
        252: log1f = 32'b01000100001111000010010011001101;
        253: log1f = 32'b01000100001111011010011000011110;
        254: log1f = 32'b01000100001111110010011101110000;
        255: log1f = 32'b01000100010000001010100011000001;
		
        
		endcase
		
    if(exp == 8'd255) begin
     if(frac == 23'd0) begin
      in_status = inf;
     end else begin
      in_status = nan;
     end
    end else if((exp == 8'd0)&&(frac == 23'd0)) begin
     in_status = zero;
    end else begin
     in_status = usual;
    end
	 
	 if(in_status == nan) begin
		 res_exp = 8'd255;
		 res_frac = {15'd0,8'd15};
		 res_sgn = 1'b0;
		 out = {res_sgn, res_exp, res_frac};
	 end else if (in_status == inf) begin
		if (sign) begin
		 res_exp = 8'd255;
       res_frac = {15'd0,8'd15};
		 res_sgn = 1'b0;
		 out = {res_sgn, res_exp, res_frac};
		end else begin
		 res_exp = 8'd255;
		 res_frac = 23'd0;
		 res_sgn = 1'b0;
		 out = {res_sgn, res_exp, res_frac};
		end
	 end else if (in_status == zero) begin
		 res_exp = 8'd255;
       res_frac = {15'd0,8'd15};
		 res_sgn = 1'b0;
		 out = {res_sgn, res_exp, res_frac};
	 end else begin
	   if (sign) begin
		  res_exp = 8'd255;
        res_frac = {15'd0,8'd15};
		  res_sgn = 1'b0;
		  out = {res_sgn, res_exp, res_frac};
		end else begin
		  out = tmp_res;
		  res_sgn= out[31];
		  res_exp = out[30:23];
		  res_frac = out[22:0];		  
		end
	 end
end


endmodule
